`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date: 2023/04/01 15:13:27
// Design Name: 
// Module Name: test_banch
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: 
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////


module test_banch();
reg clk,rstn,en;
reg [15:0] d;  
wire [15:0] m; 
MAV mav(.clk(clk),.rstn(rstn),.en(en),.d(d),.m(m));
initial begin
    d = 16'hffff;
    clk = 0;
    en = 0;
    rstn = 0;
end
always #1 clk = ~clk;
always #640000 en = ~en;

initial
begin
    #5 rstn = 1;
    #2000 d = 16'b0000_0000_0000_0010;
   #630000 d = 16'b0000_0000_0000_0010;
    #630000 d = 16'b0000_0000_0000_0011;
    #630000 d = 16'b0000_0000_0000_0011;
    #630000 d = 16'b0000_0000_0000_0101;
    #630000 d = 16'b0000_0000_0000_0010;
    #630000 d = 16'b000_0000_0000_0001;
    #630000 d = 16'b0000_0000_0000_0100;
    #630000 d = 16'b0000_0000_0000_0100;
    #630000 d = 16'b0000_0000_0000_0101;
    #630000 d = 16'b0000_0000_0000_0010;
    #630000 d = 16'b0000_0000_0000_0010;
    #630000 d = 16'b0000_0000_0000_0011;
    #630000 d = 16'b0000_0000_0000_0011;
    #630000 d = 16'b0000_0000_0000_0101;
    #630000 d = 16'b0000_0000_0000_0010;
    #630000 d = 16'b000_0000_0000_0001;
    #630000 d = 16'b0000_0000_0000_0100;
    #630000 d = 16'b0000_0000_0000_0100;
    #630000 d = 16'b0000_0000_0000_0101;
        #630000 d = 16'b0000_0000_0000_0100;
    #630000 d = 16'b0000_0000_0000_0100;
    #630000 d = 16'b0000_0000_0000_0101;
    #630000 d = 16'b0000_0000_0000_0010;
    #630000 d = 16'b0000_0000_0000_0010;
    #630000 d = 16'b0000_0000_0000_0011;
    #630000 d = 16'b0000_0000_0000_0011;
    #630000 d = 16'b0000_0000_0000_0101;
    #630000 d = 16'b0000_0000_0000_0010;
    #630000 d = 16'b000_0000_0000_0001;
    #630000 d = 16'b0000_0000_0000_0100;
    #630000 d = 16'b0000_0000_0000_0100;
    #630000 d = 16'b0000_0000_0000_0101;
end


endmodule
